module 
Dut ( 
    input [31: 0] a, 
    input clk,
    input reset, 
    output [3: 0] b 
);
endmodule
